-- Daniel Hamilton & Michael Thomas

-- SUMMARY: This testbench performs the following tests..
-- 1.) 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;